`include "cpu_types_pkg.vh"
