`ifndef CONTROL_UNIT_IF_VH
`define CONTROL_UNIT_IF_VH
